library verilog;
use verilog.vl_types.all;
entity ID_stage_sv_unit is
end ID_stage_sv_unit;
