library verilog;
use verilog.vl_types.all;
entity MDR_sv_unit is
end MDR_sv_unit;
