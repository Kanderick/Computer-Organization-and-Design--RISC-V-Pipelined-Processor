library verilog;
use verilog.vl_types.all;
entity EX_stage_sv_unit is
end EX_stage_sv_unit;
