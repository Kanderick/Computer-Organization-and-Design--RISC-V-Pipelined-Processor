library verilog;
use verilog.vl_types.all;
entity CMP_sv_unit is
end CMP_sv_unit;
