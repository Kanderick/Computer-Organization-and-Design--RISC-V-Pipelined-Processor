library verilog;
use verilog.vl_types.all;
entity mp3_cpu_sv_unit is
end mp3_cpu_sv_unit;
