library verilog;
use verilog.vl_types.all;
entity JB_hazard_detection_unit_sv_unit is
end JB_hazard_detection_unit_sv_unit;
