library verilog;
use verilog.vl_types.all;
entity control_word_reg_sv_unit is
end control_word_reg_sv_unit;
