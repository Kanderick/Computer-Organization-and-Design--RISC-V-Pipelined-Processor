library verilog;
use verilog.vl_types.all;
entity mem_access_proxy_sv_unit is
end mem_access_proxy_sv_unit;
