library verilog;
use verilog.vl_types.all;
entity control_memory_sv_unit is
end control_memory_sv_unit;
