library verilog;
use verilog.vl_types.all;
entity rdata_out_logic_sv_unit is
end rdata_out_logic_sv_unit;
