library verilog;
use verilog.vl_types.all;
entity arbitor_sv_unit is
end arbitor_sv_unit;
